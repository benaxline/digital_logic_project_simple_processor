module mov(Rx, Ry);
    input [3:0] Rx, Ry;

    

endmodule   